/*
    FULL ADDER_Module
	 
    Copyright (C) 2023  Michael Navallo Higgins

    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/

//full_adder
module f_add(a,b,carryIN,carryOUT,sum);
//declare
 input a,b,carryIN;
 output carryOUT,sum;
 wire w1,w2,w3;
 
//operation;
 h_add();



//esc
endmodule