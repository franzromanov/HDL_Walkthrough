module BCD_7(out,inp);
//start****

	//declare
	input  [3:0] inp;
	output [9:0] out;
	
//---------------------OPERATE---------------------//

//output------------------------------------------[1]
	assign out[0]=~inp[0]&~inp[1]&~inp[2]&~inp[3];

//output------------------------------------------[2]
	assign out[1]=inp[0]&~inp[1]&~inp[2]&~inp[3];

//output------------------------------------------[3]
	assign out[2]=~inp[0]&inp[1]&~inp[2]&~inp[3];

//output------------------------------------------[4]
	assign out[3]=inp[0]&inp[1]&~inp[2]&~inp[3];

//output------------------------------------------[5]
	assign out[4]=~inp[0]&~inp[1]&inp[2]&~inp[3];

//output------------------------------------------[6]
	assign out[5]=inp[0]&~inp[1]&inp[2]&~inp[3];

//output------------------------------------------[7]
	assign out[6]=~inp[0]&inp[1]&inp[2]&~inp[3];

//output------------------------------------------[8]
	assign out[7]=inp[0]&inp[1]&inp[2]&~inp[3];

//output------------------------------------------[9]
	assign out[8]=~inp[0]&~inp[1]&~inp[2]&inp[3];

//output------------------------------------------[10]
	assign out[9]=inp[0]&~inp[1]&~inp[2]&inp[3];

//-----------------------END------------------------//


//esc****
endmodule