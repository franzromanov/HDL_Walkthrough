module _OR(_OUT,A,B);
//start

 //declare
 input A,B;
 output _OUT;
 
 //operate
 assign _OUT=A|B;

//esc
endmodule