//basic_gate:NOT
module _NOT(_in,_out);
  
//declare
 input _in;
 output _out;
  
//operation
 assign _in=~_out;
  
//esc
endmodule
  
